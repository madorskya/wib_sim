library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package freq_pkg is
type t_freq is (f125, f156_25);
end package;

package body freq_pkg is

end package body;
