//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/28/2023 09:29:05 AM
// Design Name: 
// Module Name: ethernet_common_125
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ps/1ps
module ultrascale_125_gthe4_common_wrapper
(
     input  refclk,
     input  [0:0]  qpll0reset,
     output [0:0]  qpll0lock,
     output [0:0]  qpll0outclk,
     output [0:0]  qpll0outrefclk,
     input  [0:0]  qpll1reset,
     output [0:0]  qpll1lock,
     output [0:0]  qpll1outclk,
     output [0:0]  qpll1outrefclk
);

  // List of signals to connect to GT Common block

  wire [0 :0] GTHE4_COMMON_QPLL0RESET;
  wire [0 :0] GTHE4_COMMON_GTREFCLK00;
  wire [0 :0] GTHE4_COMMON_GTREFCLK01;
  wire [0 :0] GTHE4_COMMON_QPLL0LOCK;
  wire [0 :0] GTHE4_COMMON_QPLL0OUTCLK;
  wire [0 :0] GTHE4_COMMON_QPLL0OUTREFCLK;
  wire [0 :0] GTHE4_COMMON_QPLL1RESET;
  wire [0 :0] GTHE4_COMMON_QPLL1LOCK;
  wire [0 :0] GTHE4_COMMON_QPLL1OUTCLK;
  wire [0 :0] GTHE4_COMMON_QPLL1OUTREFCLK;

  // Connect only required internal signals to GT Common block
  assign GTHE4_COMMON_QPLL0RESET = qpll0reset;                  //
  assign GTHE4_COMMON_GTREFCLK00 = refclk;                      //
  assign GTHE4_COMMON_GTREFCLK01 = refclk;
  assign qpll0lock               = GTHE4_COMMON_QPLL0LOCK;      //
  assign qpll0outclk             = GTHE4_COMMON_QPLL0OUTCLK;    //
  assign qpll0outrefclk          = GTHE4_COMMON_QPLL0OUTREFCLK; // 
  assign GTHE4_COMMON_QPLL1RESET = qpll1reset;                  //
  assign qpll1lock               = GTHE4_COMMON_QPLL1LOCK;      //
  assign qpll1outclk             = GTHE4_COMMON_QPLL1OUTCLK;    //
  assign qpll1outrefclk          = GTHE4_COMMON_QPLL1OUTREFCLK; //


  xxv_ethernet_0_gt_gthe4_common_wrapper_125 xxv_ethernet_0_gt_gthe4_common_wrapper_i
  (
   .GTHE4_COMMON_BGBYPASSB(1'b1),
   .GTHE4_COMMON_BGMONITORENB(1'b1),
   .GTHE4_COMMON_BGPDB(1'b1),
   .GTHE4_COMMON_BGRCALOVRD(5'b11111),
   .GTHE4_COMMON_BGRCALOVRDENB(1'b1),
   .GTHE4_COMMON_DRPADDR(16'b0000000000000000),
   .GTHE4_COMMON_DRPCLK(1'b0),
   .GTHE4_COMMON_DRPDI(16'b0000000000000000),
   .GTHE4_COMMON_DRPDO(),
   .GTHE4_COMMON_DRPEN(1'b0),
   .GTHE4_COMMON_DRPRDY(),
   .GTHE4_COMMON_DRPWE(1'b0),
   .GTHE4_COMMON_GTGREFCLK0(1'b0),
   .GTHE4_COMMON_GTGREFCLK1(1'b0),
   .GTHE4_COMMON_GTNORTHREFCLK00(1'b0),
   .GTHE4_COMMON_GTNORTHREFCLK01(1'b0),
   .GTHE4_COMMON_GTNORTHREFCLK10(1'b0),
   .GTHE4_COMMON_GTNORTHREFCLK11(1'b0),
   .GTHE4_COMMON_GTREFCLK00(GTHE4_COMMON_GTREFCLK00),
   .GTHE4_COMMON_GTREFCLK01(1'b0),
   .GTHE4_COMMON_GTREFCLK10(1'b0),
   .GTHE4_COMMON_GTREFCLK11(1'b0),
   .GTHE4_COMMON_GTSOUTHREFCLK00(1'b0),
   .GTHE4_COMMON_GTSOUTHREFCLK01(1'b0),
   .GTHE4_COMMON_GTSOUTHREFCLK10(1'b0),
   .GTHE4_COMMON_GTSOUTHREFCLK11(1'b0),
   .GTHE4_COMMON_PCIERATEQPLL0(3'b000),
   .GTHE4_COMMON_PCIERATEQPLL1(3'b000),
   .GTHE4_COMMON_PMARSVD0(8'b00000000),
   .GTHE4_COMMON_PMARSVD1(8'b00000000),
   .GTHE4_COMMON_PMARSVDOUT0(),
   .GTHE4_COMMON_PMARSVDOUT1(),
   .GTHE4_COMMON_QPLL0CLKRSVD0(1'b0),
   .GTHE4_COMMON_QPLL0CLKRSVD1(1'b0),
   .GTHE4_COMMON_QPLL0FBCLKLOST(),
   .GTHE4_COMMON_QPLL0FBDIV(8'b00000000),
   .GTHE4_COMMON_QPLL0LOCK(GTHE4_COMMON_QPLL0LOCK),
   .GTHE4_COMMON_QPLL0LOCKDETCLK(1'b0),
   .GTHE4_COMMON_QPLL0LOCKEN(1'b1),
   .GTHE4_COMMON_QPLL0OUTCLK(GTHE4_COMMON_QPLL0OUTCLK),
   .GTHE4_COMMON_QPLL0OUTREFCLK(GTHE4_COMMON_QPLL0OUTREFCLK),
   .GTHE4_COMMON_QPLL0PD(1'b0),
   .GTHE4_COMMON_QPLL0REFCLKLOST(),
   .GTHE4_COMMON_QPLL0REFCLKSEL(3'b001),
   .GTHE4_COMMON_QPLL0RESET(GTHE4_COMMON_QPLL0RESET),
   .GTHE4_COMMON_QPLL1CLKRSVD0(1'b0),
   .GTHE4_COMMON_QPLL1CLKRSVD1(1'b0),
   .GTHE4_COMMON_QPLL1FBCLKLOST(),
   .GTHE4_COMMON_QPLL1FBDIV(8'b00000000),
   .GTHE4_COMMON_QPLL1LOCK(GTHE4_COMMON_QPLL1LOCK),
   .GTHE4_COMMON_QPLL1LOCKDETCLK(1'b0),
   .GTHE4_COMMON_QPLL1LOCKEN(1'b0),
   .GTHE4_COMMON_QPLL1OUTCLK(GTHE4_COMMON_QPLL1OUTCLK),
   .GTHE4_COMMON_QPLL1OUTREFCLK(GTHE4_COMMON_QPLL1OUTREFCLK),
   .GTHE4_COMMON_QPLL1PD(1'b1),
   .GTHE4_COMMON_QPLL1REFCLKLOST(),
   .GTHE4_COMMON_QPLL1REFCLKSEL(3'b001),
   .GTHE4_COMMON_QPLL1RESET(GTHE4_COMMON_QPLL1RESET),
   .GTHE4_COMMON_QPLLDMONITOR0(),
   .GTHE4_COMMON_QPLLDMONITOR1(),
   .GTHE4_COMMON_QPLLRSVD1(8'b00000000),
   .GTHE4_COMMON_QPLLRSVD2(5'b00000),
   .GTHE4_COMMON_QPLLRSVD3(5'b00000),
   .GTHE4_COMMON_QPLLRSVD4(8'b00000000),
   .GTHE4_COMMON_RCALENB(1'b1),
   .GTHE4_COMMON_REFCLKOUTMONITOR0(),
   .GTHE4_COMMON_REFCLKOUTMONITOR1(),
   .GTHE4_COMMON_RXRECCLK0SEL(),
   .GTHE4_COMMON_RXRECCLK1SEL(),
   .GTHE4_COMMON_SDM0DATA(25'b0100000000000000000000000),
   .GTHE4_COMMON_SDM0FINALOUT(),
   .GTHE4_COMMON_SDM0RESET(1'b0),
   .GTHE4_COMMON_SDM0TESTDATA(),
   .GTHE4_COMMON_SDM0TOGGLE(1'b0),
   .GTHE4_COMMON_SDM0WIDTH(2'b00),
   .GTHE4_COMMON_SDM1DATA(25'b0000000000000000000000000),
   .GTHE4_COMMON_SDM1FINALOUT(),
   .GTHE4_COMMON_SDM1RESET(1'b0),
   .GTHE4_COMMON_SDM1TESTDATA(),
   .GTHE4_COMMON_SDM1TOGGLE(1'b0),
   .GTHE4_COMMON_SDM1WIDTH(2'b00),
   .GTHE4_COMMON_TCONGPI(10'b0000000000),
   .GTHE4_COMMON_TCONGPO(),
   .GTHE4_COMMON_TCONPOWERUP(1'b0),
   .GTHE4_COMMON_TCONRESET(2'b00),
   .GTHE4_COMMON_TCONRSVDIN1(2'b00),
   .GTHE4_COMMON_TCONRSVDOUT0()
  );

endmodule

//ultrascale_v1_7_14_gthe4_common #(
//  .GTHE4_COMMON_AEN_QPLL0_FBDIV                 (1'b1),
//  .GTHE4_COMMON_AEN_QPLL1_FBDIV                 (1'b1),
//  .GTHE4_COMMON_AEN_SDM0TOGGLE                  (1'b0),
//  .GTHE4_COMMON_AEN_SDM1TOGGLE                  (1'b0),
//  .GTHE4_COMMON_A_SDM0TOGGLE                    (1'b0),
//  .GTHE4_COMMON_A_SDM1DATA_HIGH                 (9'b000000000),
//  .GTHE4_COMMON_A_SDM1DATA_LOW                  (16'b0000000000000000),
//  .GTHE4_COMMON_A_SDM1TOGGLE                    (1'b0),
//  .GTHE4_COMMON_BGBYPASSB_TIE_EN                (1'b0),
//  .GTHE4_COMMON_BGBYPASSB_VAL                   (1'b1),
//  .GTHE4_COMMON_BGMONITORENB_TIE_EN             (1'b0),
//  .GTHE4_COMMON_BGMONITORENB_VAL                (1'b1),
//  .GTHE4_COMMON_BGPDB_TIE_EN                    (1'b0),
//  .GTHE4_COMMON_BGPDB_VAL                       (1'b1),
//  .GTHE4_COMMON_BGRCALOVRDENB_TIE_EN            (1'b0),
//  .GTHE4_COMMON_BGRCALOVRDENB_VAL               (1'b1),
//  .GTHE4_COMMON_BGRCALOVRD_TIE_EN               (1'b0),
//  .GTHE4_COMMON_BGRCALOVRD_VAL                  (5'b11111),
//  .GTHE4_COMMON_BIAS_CFG0                       (16'b0000000000000000),
//  .GTHE4_COMMON_BIAS_CFG1                       (16'b0000000000000000),
//  .GTHE4_COMMON_BIAS_CFG2                       (16'b0000000100100100),
//  .GTHE4_COMMON_BIAS_CFG3                       (16'b0000000001000001),
//  .GTHE4_COMMON_BIAS_CFG4                       (16'b0000000000010000),
//  .GTHE4_COMMON_BIAS_CFG_RSVD                   (16'b0000000000000000),
//  .GTHE4_COMMON_COMMON_CFG0                     (16'b0000000000000000),
//  .GTHE4_COMMON_COMMON_CFG1                     (16'b0000000000000000),
//  .GTHE4_COMMON_DRPADDR_TIE_EN                  (1'b0),
//  .GTHE4_COMMON_DRPADDR_VAL                     (16'b0000000000000000),
//  .GTHE4_COMMON_DRPCLK_TIE_EN                   (1'b0),
//  .GTHE4_COMMON_DRPCLK_VAL                      (1'b0),
//  .GTHE4_COMMON_DRPDI_TIE_EN                    (1'b0),
//  .GTHE4_COMMON_DRPDI_VAL                       (16'b0000000000000000),
//  .GTHE4_COMMON_DRPEN_TIE_EN                    (1'b0),
//  .GTHE4_COMMON_DRPEN_VAL                       (1'b0),
//  .GTHE4_COMMON_DRPWE_TIE_EN                    (1'b0),
//  .GTHE4_COMMON_DRPWE_VAL                       (1'b0),
//  .GTHE4_COMMON_GTGREFCLK0_TIE_EN               (1'b0),
//  .GTHE4_COMMON_GTGREFCLK0_VAL                  (1'b0),
//  .GTHE4_COMMON_GTGREFCLK1_TIE_EN               (1'b0),
//  .GTHE4_COMMON_GTGREFCLK1_VAL                  (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK00_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK00_VAL             (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK01_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK01_VAL             (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK10_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK10_VAL             (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK11_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTNORTHREFCLK11_VAL             (1'b0),
//  .GTHE4_COMMON_GTREFCLK00_TIE_EN               (1'b0),
//  .GTHE4_COMMON_GTREFCLK00_VAL                  (1'b0),
//  .GTHE4_COMMON_GTREFCLK01_TIE_EN               (1'b0),
//  .GTHE4_COMMON_GTREFCLK01_VAL                  (1'b0),
//  .GTHE4_COMMON_GTREFCLK10_TIE_EN               (1'b0),
//  .GTHE4_COMMON_GTREFCLK10_VAL                  (1'b0),
//  .GTHE4_COMMON_GTREFCLK11_TIE_EN               (1'b0),
//  .GTHE4_COMMON_GTREFCLK11_VAL                  (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK00_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK00_VAL             (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK01_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK01_VAL             (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK10_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK10_VAL             (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK11_TIE_EN          (1'b0),
//  .GTHE4_COMMON_GTSOUTHREFCLK11_VAL             (1'b0),
//  .GTHE4_COMMON_PCIERATEQPLL0_TIE_EN            (1'b0),
//  .GTHE4_COMMON_PCIERATEQPLL0_VAL               (3'b000),
//  .GTHE4_COMMON_PCIERATEQPLL1_TIE_EN            (1'b0),
//  .GTHE4_COMMON_PCIERATEQPLL1_VAL               (3'b000),
//  .GTHE4_COMMON_PMARSVD0_TIE_EN                 (1'b0),
//  .GTHE4_COMMON_PMARSVD0_VAL                    (8'b00000000),
//  .GTHE4_COMMON_PMARSVD1_TIE_EN                 (1'b0),
//  .GTHE4_COMMON_PMARSVD1_VAL                    (8'b00000000),
//  .GTHE4_COMMON_POR_CFG                         (16'b0000000000000000),
//  .GTHE4_COMMON_PPF0_CFG                        (16'b0000011000000000),
//  .GTHE4_COMMON_PPF1_CFG                        (16'b0000011000000000),
//  .GTHE4_COMMON_QPLL0CLKOUT_RATE                ("HALF"),
//  .GTHE4_COMMON_QPLL0CLKRSVD0_TIE_EN            (1'b0),
//  .GTHE4_COMMON_QPLL0CLKRSVD0_VAL               (1'b0),
//  .GTHE4_COMMON_QPLL0CLKRSVD1_TIE_EN            (1'b0),
//  .GTHE4_COMMON_QPLL0CLKRSVD1_VAL               (1'b0),
//  .GTHE4_COMMON_QPLL0FBDIV_TIE_EN               (1'b0),
//  .GTHE4_COMMON_QPLL0FBDIV_VAL                  (8'b00000000),
//  .GTHE4_COMMON_QPLL0LOCKDETCLK_TIE_EN          (1'b0),
//  .GTHE4_COMMON_QPLL0LOCKDETCLK_VAL             (1'b0),
//  .GTHE4_COMMON_QPLL0LOCKEN_TIE_EN              (1'b0),
//  .GTHE4_COMMON_QPLL0LOCKEN_VAL                 (1'b1),
//  .GTHE4_COMMON_QPLL0PD_TIE_EN                  (1'b0),
//  .GTHE4_COMMON_QPLL0PD_VAL                     (1'b0),
//  .GTHE4_COMMON_QPLL0REFCLKSEL_TIE_EN           (1'b0),
//  .GTHE4_COMMON_QPLL0REFCLKSEL_VAL              (3'b001),
//  .GTHE4_COMMON_QPLL0RESET_TIE_EN               (1'b0),
//  .GTHE4_COMMON_QPLL0RESET_VAL                  (1'b0),
//  .GTHE4_COMMON_QPLL0_CFG0                      (16'b0011001100011100),
//  .GTHE4_COMMON_QPLL0_CFG1                      (16'b1101000000111000),
//  .GTHE4_COMMON_QPLL0_CFG1_G3                   (16'b1101000000111000),
//  .GTHE4_COMMON_QPLL0_CFG2                      (16'b0000111111000000),
//  .GTHE4_COMMON_QPLL0_CFG2_G3                   (16'b0000111111000000),
//  .GTHE4_COMMON_QPLL0_CFG3                      (16'b0000000100100000),
//  .GTHE4_COMMON_QPLL0_CFG4                      (16'b0000000000000011),
//  .GTHE4_COMMON_QPLL0_CP                        (10'b0011111111),
//  .GTHE4_COMMON_QPLL0_CP_G3                     (10'b0000001111),
//  .GTHE4_COMMON_QPLL0_FBDIV                     (66),
//  .GTHE4_COMMON_QPLL0_FBDIV_G3                  (160),
//  .GTHE4_COMMON_QPLL0_INIT_CFG0                 (16'b0000001010110010),
//  .GTHE4_COMMON_QPLL0_INIT_CFG1                 (8'b00000000),
//  .GTHE4_COMMON_QPLL0_LOCK_CFG                  (16'b0010010111101000),
//  .GTHE4_COMMON_QPLL0_LOCK_CFG_G3               (16'b0010010111101000),
//  .GTHE4_COMMON_QPLL0_LPF                       (10'b1000111111),
//  .GTHE4_COMMON_QPLL0_LPF_G3                    (10'b0111010101),
//  .GTHE4_COMMON_QPLL0_PCI_EN                    (1'b0),
//  .GTHE4_COMMON_QPLL0_RATE_SW_USE_DRP           (1'b1),
//  .GTHE4_COMMON_QPLL0_REFCLK_DIV                (1),
//  .GTHE4_COMMON_QPLL0_SDM_CFG0                  (16'b0000000010000000),
//  .GTHE4_COMMON_QPLL0_SDM_CFG1                  (16'b0000000000000000),
//  .GTHE4_COMMON_QPLL0_SDM_CFG2                  (16'b0000000000000000),
//  .GTHE4_COMMON_QPLL1CLKOUT_RATE                ("HALF"),
//  .GTHE4_COMMON_QPLL1CLKRSVD0_TIE_EN            (1'b0),
//  .GTHE4_COMMON_QPLL1CLKRSVD0_VAL               (1'b0),
//  .GTHE4_COMMON_QPLL1CLKRSVD1_TIE_EN            (1'b0),
//  .GTHE4_COMMON_QPLL1CLKRSVD1_VAL               (1'b0),
//  .GTHE4_COMMON_QPLL1FBDIV_TIE_EN               (1'b0),
//  .GTHE4_COMMON_QPLL1FBDIV_VAL                  (8'b00000000),
//  .GTHE4_COMMON_QPLL1LOCKDETCLK_TIE_EN          (1'b0),
//  .GTHE4_COMMON_QPLL1LOCKDETCLK_VAL             (1'b0),
//  .GTHE4_COMMON_QPLL1LOCKEN_TIE_EN              (1'b0),
//  .GTHE4_COMMON_QPLL1LOCKEN_VAL                 (1'b0),
//  .GTHE4_COMMON_QPLL1PD_TIE_EN                  (1'b0),
//  .GTHE4_COMMON_QPLL1PD_VAL                     (1'b1),
//  .GTHE4_COMMON_QPLL1REFCLKSEL_TIE_EN           (1'b0),
//  .GTHE4_COMMON_QPLL1REFCLKSEL_VAL              (3'b001),
//  .GTHE4_COMMON_QPLL1RESET_TIE_EN               (1'b0),
//  .GTHE4_COMMON_QPLL1RESET_VAL                  (1'b1),
//  .GTHE4_COMMON_QPLL1_CFG0                      (16'b0011001100011100),
//  .GTHE4_COMMON_QPLL1_CFG1                      (16'b1101000000111000),
//  .GTHE4_COMMON_QPLL1_CFG1_G3                   (16'b1101000000111000),
//  .GTHE4_COMMON_QPLL1_CFG2                      (16'b0000111111000011),
//  .GTHE4_COMMON_QPLL1_CFG2_G3                   (16'b0000111111000011),
//  .GTHE4_COMMON_QPLL1_CFG3                      (16'b0000000100100000),
//  .GTHE4_COMMON_QPLL1_CFG4                      (16'b0000000000000011),
//  .GTHE4_COMMON_QPLL1_CP                        (10'b0011111111),
//  .GTHE4_COMMON_QPLL1_CP_G3                     (10'b0001111111),
//  .GTHE4_COMMON_QPLL1_FBDIV                     (66),
//  .GTHE4_COMMON_QPLL1_FBDIV_G3                  (80),
//  .GTHE4_COMMON_QPLL1_INIT_CFG0                 (16'b0000001010110010),
//  .GTHE4_COMMON_QPLL1_INIT_CFG1                 (8'b00000000),
//  .GTHE4_COMMON_QPLL1_LOCK_CFG                  (16'b0010010111101000),
//  .GTHE4_COMMON_QPLL1_LOCK_CFG_G3               (16'b0010010111101000),
//  .GTHE4_COMMON_QPLL1_LPF                       (10'b1000011111),
//  .GTHE4_COMMON_QPLL1_LPF_G3                    (10'b0111010100),
//  .GTHE4_COMMON_QPLL1_PCI_EN                    (1'b0),
//  .GTHE4_COMMON_QPLL1_RATE_SW_USE_DRP           (1'b1),
//  .GTHE4_COMMON_QPLL1_REFCLK_DIV                (1),
//  .GTHE4_COMMON_QPLL1_SDM_CFG0                  (16'b0000000010000000),
//  .GTHE4_COMMON_QPLL1_SDM_CFG1                  (16'b0000000000000000),
//  .GTHE4_COMMON_QPLL1_SDM_CFG2                  (16'b0000000000000000),
//  .GTHE4_COMMON_QPLLRSVD1_TIE_EN                (1'b0),
//  .GTHE4_COMMON_QPLLRSVD1_VAL                   (8'b00000000),
//  .GTHE4_COMMON_QPLLRSVD2_TIE_EN                (1'b0),
//  .GTHE4_COMMON_QPLLRSVD2_VAL                   (5'b00000),
//  .GTHE4_COMMON_QPLLRSVD3_TIE_EN                (1'b0),
//  .GTHE4_COMMON_QPLLRSVD3_VAL                   (5'b00000),
//  .GTHE4_COMMON_QPLLRSVD4_TIE_EN                (1'b0),
//  .GTHE4_COMMON_QPLLRSVD4_VAL                   (8'b00000000),
//  .GTHE4_COMMON_RCALENB_TIE_EN                  (1'b0),
//  .GTHE4_COMMON_RCALENB_VAL                     (1'b1),
//  .GTHE4_COMMON_RSVD_ATTR0                      (16'b0000000000000000),
//  .GTHE4_COMMON_RSVD_ATTR1                      (16'b0000000000000000),
//  .GTHE4_COMMON_RSVD_ATTR2                      (16'b0000000000000000),
//  .GTHE4_COMMON_RSVD_ATTR3                      (16'b0000000000000000),
//  .GTHE4_COMMON_RXRECCLKOUT0_SEL                (2'b00),
//  .GTHE4_COMMON_RXRECCLKOUT1_SEL                (2'b00),
//  .GTHE4_COMMON_SARC_ENB                        (1'b0),
//  .GTHE4_COMMON_SARC_SEL                        (1'b0),
//  .GTHE4_COMMON_SDM0DATA_TIE_EN                 (1'b0),
//  .GTHE4_COMMON_SDM0DATA_VAL                    (25'b0000000000000000000000000),
//  .GTHE4_COMMON_SDM0INITSEED0_0                 (16'b0000000100010001),
//  .GTHE4_COMMON_SDM0INITSEED0_1                 (9'b000010001),
//  .GTHE4_COMMON_SDM0RESET_TIE_EN                (1'b0),
//  .GTHE4_COMMON_SDM0RESET_VAL                   (1'b0),
//  .GTHE4_COMMON_SDM0TOGGLE_TIE_EN               (1'b0),
//  .GTHE4_COMMON_SDM0TOGGLE_VAL                  (1'b0),
//  .GTHE4_COMMON_SDM0WIDTH_TIE_EN                (1'b0),
//  .GTHE4_COMMON_SDM0WIDTH_VAL                   (2'b00),
//  .GTHE4_COMMON_SDM1DATA_TIE_EN                 (1'b0),
//  .GTHE4_COMMON_SDM1DATA_VAL                    (25'b0000000000000000000000000),
//  .GTHE4_COMMON_SDM1INITSEED0_0                 (16'b0000000100010001),
//  .GTHE4_COMMON_SDM1INITSEED0_1                 (9'b000010001),
//  .GTHE4_COMMON_SDM1RESET_TIE_EN                (1'b0),
//  .GTHE4_COMMON_SDM1RESET_VAL                   (1'b0),
//  .GTHE4_COMMON_SDM1TOGGLE_TIE_EN               (1'b0),
//  .GTHE4_COMMON_SDM1TOGGLE_VAL                  (1'b0),
//  .GTHE4_COMMON_SDM1WIDTH_TIE_EN                (1'b0),
//  .GTHE4_COMMON_SDM1WIDTH_VAL                   (2'b00),
//  .GTHE4_COMMON_SIM_DEVICE                      ("ULTRASCALE_PLUS"),
//  .GTHE4_COMMON_SIM_MODE                        ("FAST"),
//  .GTHE4_COMMON_SIM_RESET_SPEEDUP               ("TRUE"),
//  .GTHE4_COMMON_TCONGPI_TIE_EN                  (1'b0),
//  .GTHE4_COMMON_TCONGPI_VAL                     (10'b0000000000),
//  .GTHE4_COMMON_TCONPOWERUP_TIE_EN              (1'b0),
//  .GTHE4_COMMON_TCONPOWERUP_VAL                 (1'b0),
//  .GTHE4_COMMON_TCONRESET_TIE_EN                (1'b0),
//  .GTHE4_COMMON_TCONRESET_VAL                   (2'b00),
//  .GTHE4_COMMON_TCONRSVDIN1_TIE_EN              (1'b0),
//  .GTHE4_COMMON_TCONRSVDIN1_VAL                 (2'b00)
//) common_inst (

//  // inputs
//        .GTHE4_COMMON_BGBYPASSB         (1'b1),
//        .GTHE4_COMMON_BGMONITORENB      (1'b1),
//        .GTHE4_COMMON_BGPDB             (1'b1),
//        .GTHE4_COMMON_BGRCALOVRD        (5'b11111),
//        .GTHE4_COMMON_BGRCALOVRDENB     (1'b1),
//        .GTHE4_COMMON_DRPADDR           (16'b0000000000000000),
//        .GTHE4_COMMON_DRPCLK            (1'b0),
//        .GTHE4_COMMON_DRPDI             (16'b0000000000000000),
//        .GTHE4_COMMON_DRPEN             (1'b0),
//        .GTHE4_COMMON_DRPWE             (1'b0),
//        .GTHE4_COMMON_GTGREFCLK0        (1'b0),
//        .GTHE4_COMMON_GTGREFCLK1        (1'b0),
//        .GTHE4_COMMON_GTNORTHREFCLK00   (1'b0),
//        .GTHE4_COMMON_GTNORTHREFCLK01   (1'b0),
//        .GTHE4_COMMON_GTNORTHREFCLK10   (1'b0),
//        .GTHE4_COMMON_GTNORTHREFCLK11   (1'b0),
//        .GTHE4_COMMON_GTREFCLK00        (GTHE4_COMMON_GTREFCLK00),
//        .GTHE4_COMMON_GTREFCLK01        (1'b0),
//        .GTHE4_COMMON_GTREFCLK10        (1'b0),
//        .GTHE4_COMMON_GTREFCLK11        (1'b0),
//        .GTHE4_COMMON_GTSOUTHREFCLK00   (1'b0),
//        .GTHE4_COMMON_GTSOUTHREFCLK01   (1'b0),
//        .GTHE4_COMMON_GTSOUTHREFCLK10   (1'b0),
//        .GTHE4_COMMON_GTSOUTHREFCLK11   (1'b0),
//        .GTHE4_COMMON_PCIERATEQPLL0     (3'b000),
//        .GTHE4_COMMON_PCIERATEQPLL1     (3'b000),
//        .GTHE4_COMMON_PMARSVD0          (8'b00000000),
//        .GTHE4_COMMON_PMARSVD1          (8'b00000000),
//        .GTHE4_COMMON_QPLL0CLKRSVD0     (1'b0),
//        .GTHE4_COMMON_QPLL0CLKRSVD1     (1'b0),
//        .GTHE4_COMMON_QPLL0FBDIV        (8'b00000000),
//        .GTHE4_COMMON_QPLL0LOCKDETCLK   (1'b0),
//        .GTHE4_COMMON_QPLL0LOCKEN       (1'b1),
//        .GTHE4_COMMON_QPLL0PD           (1'b0),
//        .GTHE4_COMMON_QPLL0REFCLKSEL    (3'b001),
//        .GTHE4_COMMON_QPLL0RESET        (GTHE4_COMMON_QPLL0RESET),
//        .GTHE4_COMMON_QPLL1CLKRSVD0     (1'b0),
//        .GTHE4_COMMON_QPLL1CLKRSVD1     (1'b0),
//        .GTHE4_COMMON_QPLL1FBDIV        (8'b00000000),
//        .GTHE4_COMMON_QPLL1LOCKDETCLK   (1'b0),
//        .GTHE4_COMMON_QPLL1LOCKEN       (1'b0),
//        .GTHE4_COMMON_QPLL1PD           (1'b1),
//        .GTHE4_COMMON_QPLL1REFCLKSEL    (3'b001),
//        .GTHE4_COMMON_QPLL1RESET        (GTHE4_COMMON_QPLL1RESET),
//        .GTHE4_COMMON_QPLLRSVD1         (8'b00000000),
//        .GTHE4_COMMON_QPLLRSVD2         (5'b00000),
//        .GTHE4_COMMON_QPLLRSVD3         (5'b00000),
//        .GTHE4_COMMON_QPLLRSVD4         (8'b00000000),
//        .GTHE4_COMMON_RCALENB           (1'b1),
//        .GTHE4_COMMON_SDM0DATA          (25'b0000000000000000000000000),
//        .GTHE4_COMMON_SDM0RESET         (1'b0),
//        .GTHE4_COMMON_SDM0TOGGLE        (1'b0),
//        .GTHE4_COMMON_SDM0WIDTH         (2'b00),
//        .GTHE4_COMMON_SDM1DATA          (25'b0000000000000000000000000),
//        .GTHE4_COMMON_SDM1RESET         (1'b0),
//        .GTHE4_COMMON_SDM1TOGGLE        (1'b0),
//        .GTHE4_COMMON_SDM1WIDTH         (2'b00),
//        .GTHE4_COMMON_TCONGPI           (10'b0000000000),
//        .GTHE4_COMMON_TCONPOWERUP       (1'b0),
//        .GTHE4_COMMON_TCONRESET         (2'b00),
//        .GTHE4_COMMON_TCONRSVDIN1       (2'b00),
//  // outputs
//        .GTHE4_COMMON_DRPDO             (),
//        .GTHE4_COMMON_DRPRDY            (),
//        .GTHE4_COMMON_PMARSVDOUT0       (),
//        .GTHE4_COMMON_PMARSVDOUT1       (),
//        .GTHE4_COMMON_QPLL0FBCLKLOST    (),
//        .GTHE4_COMMON_QPLL0LOCK         (GTHE4_COMMON_QPLL0LOCK),     
//        .GTHE4_COMMON_QPLL0OUTCLK       (GTHE4_COMMON_QPLL0OUTCLK),   
//        .GTHE4_COMMON_QPLL0OUTREFCLK    (GTHE4_COMMON_QPLL0OUTREFCLK),
//        .GTHE4_COMMON_QPLL0REFCLKLOST   (),
//        .GTHE4_COMMON_QPLL1FBCLKLOST    (),
//        .GTHE4_COMMON_QPLL1LOCK         (GTHE4_COMMON_QPLL1LOCK),     
//        .GTHE4_COMMON_QPLL1OUTCLK       (GTHE4_COMMON_QPLL1OUTCLK),   
//        .GTHE4_COMMON_QPLL1OUTREFCLK    (GTHE4_COMMON_QPLL1OUTREFCLK),
//        .GTHE4_COMMON_QPLL1REFCLKLOST   (),
//        .GTHE4_COMMON_QPLLDMONITOR0     (),
//        .GTHE4_COMMON_QPLLDMONITOR1     (),
//        .GTHE4_COMMON_REFCLKOUTMONITOR0 (),
//        .GTHE4_COMMON_REFCLKOUTMONITOR1 (),
//        .GTHE4_COMMON_RXRECCLK0SEL      (),
//        .GTHE4_COMMON_RXRECCLK1SEL      (),
//        .GTHE4_COMMON_SDM0FINALOUT      (),
//        .GTHE4_COMMON_SDM0TESTDATA      (),
//        .GTHE4_COMMON_SDM1FINALOUT      (),
//        .GTHE4_COMMON_SDM1TESTDATA      (),
//        .GTHE4_COMMON_TCONGPO           (),
//        .GTHE4_COMMON_TCONRSVDOUT0      ()
//);
