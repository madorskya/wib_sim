
// file: wib_ibert_coldata.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_wib_ibert_coldata
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_wib_ibert_coldata
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////

`define C_NUM_GTH_QUADS 4
`define C_GTH_REFCLKS_USED 4
module example_wib_ibert_coldata
(
  // GT top level ports
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txn_o,
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txp_o,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]    	gth_rxn_i,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]   	gth_rxp_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0n_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1n_i
);

  //
  // Ibert refclk internal signals
  //
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk1_i;        	
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk11_i; 
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk1_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_1_i;
  wire                        gth_sysclk_i;


  //
  // Refclk IBUFDS instantiations
  //
    IBUFDS_GTE4 u_buf_gth_q3_clk0
      (
        .O            (gth_refclk0_i[0]),
        .ODIV2        (gth_odiv2_0_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[0]),
        .IB           (gth_refclk0n_i[0])
      );

    IBUFDS_GTE4 u_buf_gth_q3_clk1
      (
        .O            (gth_refclk1_i[0]),
        .ODIV2        (gth_odiv2_1_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[0]),
        .IB           (gth_refclk1n_i[0])
      );
    IBUFDS_GTE4 u_buf_gth_q5_clk0
      (
        .O            (gth_refclk0_i[1]),
        .ODIV2        (gth_odiv2_0_i[1]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[1]),
        .IB           (gth_refclk0n_i[1])
      );

    IBUFDS_GTE4 u_buf_gth_q5_clk1
      (
        .O            (gth_refclk1_i[1]),
        .ODIV2        (gth_odiv2_1_i[1]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[1]),
        .IB           (gth_refclk1n_i[1])
      );
    IBUFDS_GTE4 u_buf_gth_q6_clk0
      (
        .O            (gth_refclk0_i[2]),
        .ODIV2        (gth_odiv2_0_i[2]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[2]),
        .IB           (gth_refclk0n_i[2])
      );

    IBUFDS_GTE4 u_buf_gth_q6_clk1
      (
        .O            (gth_refclk1_i[2]),
        .ODIV2        (gth_odiv2_1_i[2]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[2]),
        .IB           (gth_refclk1n_i[2])
      );
    IBUFDS_GTE4 u_buf_gth_q7_clk0
      (
        .O            (gth_refclk0_i[3]),
        .ODIV2        (gth_odiv2_0_i[3]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[3]),
        .IB           (gth_refclk0n_i[3])
      );

    IBUFDS_GTE4 u_buf_gth_q7_clk1
      (
        .O            (gth_refclk1_i[3]),
        .ODIV2        (gth_odiv2_1_i[3]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[3]),
        .IB           (gth_refclk1n_i[3])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gth_qrefclk0_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk1_i[0] = gth_refclk1_i[0];
  assign gth_qnorthrefclk0_i[0] = 1'b0;
  assign gth_qnorthrefclk1_i[0] = 1'b0;
  assign gth_qsouthrefclk0_i[0] = 1'b0;
  assign gth_qsouthrefclk1_i[0] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk10_i[0] = gth_refclk1_i[0];
  assign gth_qrefclk01_i[0] = 1'b0;
  assign gth_qrefclk11_i[0] = 1'b0;  
  assign gth_qnorthrefclk00_i[0] = 1'b0;
  assign gth_qnorthrefclk10_i[0] = 1'b0;
  assign gth_qnorthrefclk01_i[0] = 1'b0;
  assign gth_qnorthrefclk11_i[0] = 1'b0;  
  assign gth_qsouthrefclk00_i[0] = 1'b0;
  assign gth_qsouthrefclk10_i[0] = 1'b0;  
  assign gth_qsouthrefclk01_i[0] = 1'b0;
  assign gth_qsouthrefclk11_i[0] = 1'b0; 
 

  assign gth_qrefclk0_i[1] = gth_refclk0_i[1];
  assign gth_qrefclk1_i[1] = gth_refclk1_i[1];
  assign gth_qnorthrefclk0_i[1] = 1'b0;
  assign gth_qnorthrefclk1_i[1] = 1'b0;
  assign gth_qsouthrefclk0_i[1] = 1'b0;
  assign gth_qsouthrefclk1_i[1] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[1] = gth_refclk0_i[1];
  assign gth_qrefclk10_i[1] = gth_refclk1_i[1];
  assign gth_qrefclk01_i[1] = 1'b0;
  assign gth_qrefclk11_i[1] = 1'b0;  
  assign gth_qnorthrefclk00_i[1] = 1'b0;
  assign gth_qnorthrefclk10_i[1] = 1'b0;
  assign gth_qnorthrefclk01_i[1] = 1'b0;
  assign gth_qnorthrefclk11_i[1] = 1'b0;  
  assign gth_qsouthrefclk00_i[1] = 1'b0;
  assign gth_qsouthrefclk10_i[1] = 1'b0;  
  assign gth_qsouthrefclk01_i[1] = 1'b0;
  assign gth_qsouthrefclk11_i[1] = 1'b0; 
 

  assign gth_qrefclk0_i[2] = gth_refclk0_i[2];
  assign gth_qrefclk1_i[2] = gth_refclk1_i[2];
  assign gth_qnorthrefclk0_i[2] = 1'b0;
  assign gth_qnorthrefclk1_i[2] = 1'b0;
  assign gth_qsouthrefclk0_i[2] = 1'b0;
  assign gth_qsouthrefclk1_i[2] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[2] = gth_refclk0_i[2];
  assign gth_qrefclk10_i[2] = gth_refclk1_i[2];
  assign gth_qrefclk01_i[2] = 1'b0;
  assign gth_qrefclk11_i[2] = 1'b0;  
  assign gth_qnorthrefclk00_i[2] = 1'b0;
  assign gth_qnorthrefclk10_i[2] = 1'b0;
  assign gth_qnorthrefclk01_i[2] = 1'b0;
  assign gth_qnorthrefclk11_i[2] = 1'b0;  
  assign gth_qsouthrefclk00_i[2] = 1'b0;
  assign gth_qsouthrefclk10_i[2] = 1'b0;  
  assign gth_qsouthrefclk01_i[2] = 1'b0;
  assign gth_qsouthrefclk11_i[2] = 1'b0; 
 

  assign gth_qrefclk0_i[3] = gth_refclk0_i[3];
  assign gth_qrefclk1_i[3] = gth_refclk1_i[3];
  assign gth_qnorthrefclk0_i[3] = 1'b0;
  assign gth_qnorthrefclk1_i[3] = 1'b0;
  assign gth_qsouthrefclk0_i[3] = 1'b0;
  assign gth_qsouthrefclk1_i[3] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[3] = gth_refclk0_i[3];
  assign gth_qrefclk10_i[3] = gth_refclk1_i[3];
  assign gth_qrefclk01_i[3] = 1'b0;
  assign gth_qrefclk11_i[3] = 1'b0;  
  assign gth_qnorthrefclk00_i[3] = 1'b0;
  assign gth_qnorthrefclk10_i[3] = 1'b0;
  assign gth_qnorthrefclk01_i[3] = 1'b0;
  assign gth_qnorthrefclk11_i[3] = 1'b0;  
  assign gth_qsouthrefclk00_i[3] = 1'b0;
  assign gth_qsouthrefclk10_i[3] = 1'b0;  
  assign gth_qsouthrefclk01_i[3] = 1'b0;
  assign gth_qsouthrefclk11_i[3] = 1'b0; 
 

    BUFG_GT u_gth_sysclk_internal
      (
        .I        (gth_odiv2_0_i[0]),
        .O        (gth_sysclk_i),
        .CE       (1'b1),
        .CEMASK   (1'b0),
        .CLR      (1'b0),
        .CLRMASK  (1'b0),
        .DIV      (3'b000)
      );


  //
  // IBERT core instantiation
  //
  wib_ibert_coldata u_ibert_gth_core
    (
      .txn_o(gth_txn_o),
      .txp_o(gth_txp_o),
      .rxn_i(gth_rxn_i),
      .rxp_i(gth_rxp_i),
      .clk(gth_sysclk_i),
      .gtrefclk0_i(gth_qrefclk0_i),
      .gtrefclk1_i(gth_qrefclk1_i),
      .gtnorthrefclk0_i(gth_qnorthrefclk0_i),
      .gtnorthrefclk1_i(gth_qnorthrefclk1_i),
      .gtsouthrefclk0_i(gth_qsouthrefclk0_i),
      .gtsouthrefclk1_i(gth_qsouthrefclk1_i),
      .gtrefclk00_i(gth_qrefclk00_i),
      .gtrefclk10_i(gth_qrefclk10_i),
      .gtrefclk01_i(gth_qrefclk01_i),
      .gtrefclk11_i(gth_qrefclk11_i),
      .gtnorthrefclk00_i(gth_qnorthrefclk00_i),
      .gtnorthrefclk10_i(gth_qnorthrefclk10_i),
      .gtnorthrefclk01_i(gth_qnorthrefclk01_i),
      .gtnorthrefclk11_i(gth_qnorthrefclk11_i),
      .gtsouthrefclk00_i(gth_qsouthrefclk00_i),
      .gtsouthrefclk10_i(gth_qsouthrefclk10_i),
      .gtsouthrefclk01_i(gth_qsouthrefclk01_i),
      .gtsouthrefclk11_i(gth_qsouthrefclk11_i)
    );

endmodule
